library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
--use IEEE.MATH_REAL.ALL  ;
entity UART_RX is
  generic(
    SYSTEM_SPEED : integer := 4; --50e6;   	-- clock speed, in Hz 	--for simmulation setting = 4
    BAUDRATE     : integer := 1);--9600 	   -- baudrate 				--for simmulation setting = 1
  port(
    clk_i   : in  std_logic;	-- system clock 							
    rst_i   : in  std_logic;	-- synchronous reset, active-high
    req_o   : out std_logic := '0'; 	-- Rx req
    data_o  : out std_logic_vector(7 downto 0); -- Rx data
	 sampling_rx : out std_logic := '0'; 
    rx      : in std_logic );	-- Rx input
end UART_RX;
architecture behave of UART_RX is
  constant MAX_COUNTER: integer := (SYSTEM_SPEED / BAUDRATE);
   type state_type is (
     WAIT_FOR_RX_START, 
     WAIT_HALF_BIT,
     RECEIVE_BITS,
     WAIT_FOR_STOP_BIT );

  signal state : state_type := WAIT_FOR_RX_START;
  signal baudrate_counter  : integer range 0 to max_counter := 0;
  signal bit_counter : integer range 0 to 7 := 0;
  signal receive_register : std_logic_vector(7 downto 0) := (others => '0');

begin
  process (clk_i)
  begin
    if rising_edge(clk_i) then
      if rst_i = '0' then
        state  <= WAIT_FOR_RX_START;
        data_o <= (others => '0');
        req_o  <= '0';
      else
        case state is
		  
          when WAIT_FOR_RX_START =>
            if rx = '0' then
              -- start bit received, wait for a half bit time
              -- to sample bits in the middle of the signal
              state <= WAIT_HALF_BIT;
              baudrate_counter <= (MAX_COUNTER / 2) - 1;
				  req_o  <= '1';
            end if;
				
          when WAIT_HALF_BIT =>
            if baudrate_counter = 0 then
              -- now we are in the middle of the start bit,
              -- wait a full bit for the middle of the first bit
              state <= RECEIVE_BITS;
              bit_counter <= 7;
              baudrate_counter <= MAX_COUNTER - 1;
            else
              baudrate_counter <= baudrate_counter - 1;
            end if;
				
          when RECEIVE_BITS =>
            -- sample a bit
            if baudrate_counter = 0 then
              receive_register <= rx & receive_register(7 downto 1); --shift right sequence for keep lsb first
				   sampling_rx <= '1';
              if bit_counter = 0 then
                state <= WAIT_FOR_STOP_BIT;
              else
                bit_counter <= bit_counter - 1;
              end if;
              baudrate_counter <= MAX_COUNTER - 1;
            else
              baudrate_counter <= baudrate_counter - 1;
				  sampling_rx <= '0';
            end if;
            
          when WAIT_FOR_STOP_BIT =>
            -- wait for stop bit
            if baudrate_counter = 0 then
              if rx = '1' then
                data_o <= receive_register;
                req_o  <= '0';
					 state <= WAIT_FOR_RX_START;
              end if;  
            else
              baudrate_counter <= baudrate_counter - 1;
            end if;
        end case;
      end if;
    end if;
  end process;

end behave;