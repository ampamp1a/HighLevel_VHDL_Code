--VGAPLL_inst : VGAPLL PORT MAP (
--		areset	 => areset_sig,
--		inclk0	 => inclk0_sig,
--		c0	 => c0_sig
--	);
